`define SERIAL
`undef SERIAL
